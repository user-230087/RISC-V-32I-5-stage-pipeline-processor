module Adder(input [31:0] A,B,
output [31:0] op
    );
    assign op = A + B;
endmodule